module PMESH_L2_ILA__DOT__STORE_REQ(
__START__,
clk,
msg1_data,
msg1_source,
msg1_tag,
msg1_type,
msg1_valid,
msg2_ready,
msg3_data,
msg3_source,
msg3_tag,
msg3_type,
msg3_valid,
nondet___unknown__1_n78,
rst,
__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__,
__ILA_PMESH_L2_ILA_valid__,
msg1_ready,
msg3_ready,
msg2_type,
msg2_valid,
cache_tag,
cache_vd,
cache_state,
cache_data,
cache_owner,
share_list,
cur_msg_state,
cur_msg_type,
cur_msg_source,
cur_msg_tag,
__COUNTER_start__n15
);
input            __START__;
input            clk;
input     [63:0] msg1_data;
input      [5:0] msg1_source;
input     [25:0] msg1_tag;
input      [7:0] msg1_type;
input            msg1_valid;
input            msg2_ready;
input     [63:0] msg3_data;
input      [5:0] msg3_source;
input     [25:0] msg3_tag;
input      [7:0] msg3_type;
input            msg3_valid;
input      [5:0] nondet___unknown__1_n78;
input            rst;
output            __ILA_PMESH_L2_ILA_decode_of_STORE_REQ__;
output            __ILA_PMESH_L2_ILA_valid__;
output reg            msg1_ready;
output reg            msg3_ready;
output reg      [7:0] msg2_type;
output reg            msg2_valid;
output reg     [25:0] cache_tag;
output reg      [1:0] cache_vd;
output reg      [1:0] cache_state;
output reg     [63:0] cache_data;
output reg      [5:0] cache_owner;
output reg     [63:0] share_list;
output reg      [1:0] cur_msg_state;
output reg      [7:0] cur_msg_type;
output reg      [5:0] cur_msg_source;
output reg     [25:0] cur_msg_tag;
output reg      [7:0] __COUNTER_start__n15;
wire            __ILA_PMESH_L2_ILA_decode_of_STORE_REQ__;
wire            __ILA_PMESH_L2_ILA_valid__;
wire            __START__;
wire            bv_1_1_n0__$303;
wire      [1:0] bv_2_0_n6__$59;
wire      [1:0] bv_2_1_n31__$97;
wire      [1:0] bv_2_2_n10__$63;
wire      [1:0] bv_2_3_n21__$105;
wire      [7:0] bv_8_17_n34__$75;
wire      [7:0] bv_8_18_n33__$77;
wire      [7:0] bv_8_19_n29__$79;
wire      [7:0] bv_8_20_n28__$81;
wire      [7:0] bv_8_29_n43__$93;
wire      [7:0] bv_8_2_n4__$65;
(* keep *) wire     [63:0] cache_data_randinit;
(* keep *) wire      [5:0] cache_owner_randinit;
(* keep *) wire      [1:0] cache_state_randinit;
(* keep *) wire     [25:0] cache_tag_randinit;
(* keep *) wire      [1:0] cache_vd_randinit;
wire            clk;
(* keep *) wire      [5:0] cur_msg_source_randinit;
(* keep *) wire      [1:0] cur_msg_state_randinit;
(* keep *) wire     [25:0] cur_msg_tag_randinit;
(* keep *) wire      [7:0] cur_msg_type_randinit;
wire     [63:0] msg1_data;
(* keep *) wire            msg1_ready_randinit;
wire      [5:0] msg1_source;
wire     [25:0] msg1_tag;
wire      [7:0] msg1_type;
wire            msg1_valid;
wire            msg2_ready;
(* keep *) wire      [7:0] msg2_type_randinit;
(* keep *) wire            msg2_valid_randinit;
wire     [63:0] msg3_data;
(* keep *) wire            msg3_ready_randinit;
wire      [5:0] msg3_source;
wire     [25:0] msg3_tag;
wire      [7:0] msg3_type;
wire            msg3_valid;
wire            n11__$319;
wire            n12__$321;
wire            n13__$322;
wire            n14__$323;
wire            n16__$137;
wire     [25:0] n17__$139;
wire            n18__$140;
wire            n19__$142;
wire            n1__$305;
wire            n20__$143;
wire            n22__$145;
wire            n23__$147;
wire            n24__$148;
wire            n25__$396;
wire            n26__$398;
wire            n27__$400;
wire            n2__$309;
wire      [7:0] n30__$402;
wire            n32__$403;
wire      [7:0] n35__$405;
wire      [7:0] n36__$406;
wire            n37__$149;
wire            n38__$409;
wire            n39__$411;
wire            n3__$311;
wire            n40__$121;
wire      [5:0] n41__$123;
wire            n42__$124;
wire      [7:0] n44__$413;
wire            n45__$414;
wire      [7:0] n46__$416;
wire      [7:0] n47__$417;
wire      [7:0] n48__$418;
wire      [7:0] n49__$419;
wire            n50__$360;
wire            n51__$362;
wire      [1:0] n52__$364;
wire      [1:0] n53__$365;
wire            n54__$126;
wire     [25:0] n55__$128;
wire            n56__$129;
wire            n57__$131;
wire            n58__$133;
wire            n59__$135;
wire            n5__$312;
wire            n60__$136;
wire            n61__$352;
wire            n62__$354;
wire      [1:0] n63__$356;
wire      [1:0] n64__$357;
wire            n65__$326;
wire            n66__$328;
wire            n67__$330;
wire            n68__$331;
wire            n69__$332;
wire            n70__$333;
wire            n71__$335;
wire            n72__$336;
wire            n73__$366;
wire            n74__$368;
wire      [5:0] n75__$370;
wire      [5:0] n76__$371;
wire            n77__$372;
wire      [5:0] n79__$376;
wire            n7__$314;
wire      [5:0] n80__$392;
wire      [5:0] n81__$393;
wire      [1:0] n82__$349;
wire            n83__$337;
wire            n84__$339;
wire      [7:0] n85__$340;
wire            n86__$345;
wire            n87__$347;
wire      [5:0] n88__$348;
wire            n89__$341;
wire            n8__$316;
wire            n90__$343;
wire     [25:0] n91__$344;
wire            n9__$317;
wire      [5:0] nondet___unknown__1_n78;
wire            rst;
(* keep *) wire     [63:0] share_list_randinit;
assign __ILA_PMESH_L2_ILA_valid__ = 1'b1 ;
assign bv_1_1_n0__$303 = 1'h1 ;
assign n1__$305 =  ( msg1_ready ) == ( bv_1_1_n0__$303 )  ;
assign n2__$309 =  ( msg1_valid ) == ( bv_1_1_n0__$303 )  ;
assign n3__$311 =  ( n1__$305 ) & (n2__$309 )  ;
assign bv_8_2_n4__$65 = 8'h2 ;
assign n5__$312 =  ( msg1_type ) == ( bv_8_2_n4__$65 )  ;
assign bv_2_0_n6__$59 = 2'h0 ;
assign n7__$314 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n8__$316 =  ( n5__$312 ) & (n7__$314 )  ;
assign n9__$317 =  ( cur_msg_type ) == ( bv_8_2_n4__$65 )  ;
assign bv_2_2_n10__$63 = 2'h2 ;
assign n11__$319 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n12__$321 =  ( n9__$317 ) & (n11__$319 )  ;
assign n13__$322 =  ( n8__$316 ) | ( n12__$321 )  ;
assign n14__$323 =  ( n3__$311 ) & (n13__$322 )  ;
assign __ILA_PMESH_L2_ILA_decode_of_STORE_REQ__ = n14__$323 ;
assign n16__$137 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n17__$139 =  ( n16__$137 ) ? ( msg1_tag ) : ( cur_msg_tag ) ;
assign n18__$140 =  ( n17__$139 ) == ( cache_tag )  ;
assign n19__$142 = ~ ( n18__$140 )  ;
assign n20__$143 =  ( cache_vd ) == ( bv_2_2_n10__$63 )  ;
assign bv_2_3_n21__$105 = 2'h3 ;
assign n22__$145 =  ( cache_vd ) == ( bv_2_3_n21__$105 )  ;
assign n23__$147 =  ( n20__$143 ) | ( n22__$145 )  ;
assign n24__$148 =  ( n19__$142 ) & (n23__$147 )  ;
assign n25__$396 =  ( n24__$148 ) == ( 1'b1 )  ;
assign n26__$398 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n27__$400 =  ( cache_vd ) == ( bv_2_3_n21__$105 )  ;
assign bv_8_20_n28__$81 = 8'h14 ;
assign bv_8_19_n29__$79 = 8'h13 ;
assign n30__$402 =  ( n27__$400 ) ? ( bv_8_20_n28__$81 ) : ( bv_8_19_n29__$79 ) ;
assign bv_2_1_n31__$97 = 2'h1 ;
assign n32__$403 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign bv_8_18_n33__$77 = 8'h12 ;
assign bv_8_17_n34__$75 = 8'h11 ;
assign n35__$405 =  ( n32__$403 ) ? ( bv_8_18_n33__$77 ) : ( bv_8_17_n34__$75 ) ;
assign n36__$406 =  ( n26__$398 ) ? ( n30__$402 ) : ( n35__$405 ) ;
assign n37__$149 =  ( cache_vd ) == ( bv_2_0_n6__$59 )  ;
assign n38__$409 =  ( n37__$149 ) == ( 1'b1 )  ;
assign n39__$411 =  ( cache_state ) == ( bv_2_2_n10__$63 )  ;
assign n40__$121 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n41__$123 =  ( n40__$121 ) ? ( msg1_source ) : ( cur_msg_source ) ;
assign n42__$124 =  ( n41__$123 ) == ( cache_owner )  ;
assign bv_8_29_n43__$93 = 8'h1d ;
assign n44__$413 =  ( n42__$124 ) ? ( bv_8_29_n43__$93 ) : ( bv_8_17_n34__$75 ) ;
assign n45__$414 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign n46__$416 =  ( n45__$414 ) ? ( bv_8_18_n33__$77 ) : ( bv_8_29_n43__$93 ) ;
assign n47__$417 =  ( n39__$411 ) ? ( n44__$413 ) : ( n46__$416 ) ;
assign n48__$418 =  ( n38__$409 ) ? ( bv_8_19_n29__$79 ) : ( n47__$417 ) ;
assign n49__$419 =  ( n25__$396 ) ? ( n36__$406 ) : ( n48__$418 ) ;
assign n50__$360 =  ( n24__$148 ) == ( 1'b1 )  ;
assign n51__$362 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n52__$364 =  ( n51__$362 ) ? ( bv_2_0_n6__$59 ) : ( cache_vd ) ;
assign n53__$365 =  ( n50__$360 ) ? ( n52__$364 ) : ( cache_vd ) ;
assign n54__$126 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n55__$128 =  ( n54__$126 ) ? ( msg1_tag ) : ( cur_msg_tag ) ;
assign n56__$129 =  ( n55__$128 ) == ( cache_tag )  ;
assign n57__$131 =  ( cache_vd ) == ( bv_2_2_n10__$63 )  ;
assign n58__$133 =  ( cache_vd ) == ( bv_2_3_n21__$105 )  ;
assign n59__$135 =  ( n57__$131 ) | ( n58__$133 )  ;
assign n60__$136 =  ( n56__$129 ) & (n59__$135 )  ;
assign n61__$352 =  ( n60__$136 ) == ( 1'b1 )  ;
assign n62__$354 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n63__$356 =  ( n62__$354 ) ? ( bv_2_2_n10__$63 ) : ( cache_state ) ;
assign n64__$357 =  ( n61__$352 ) ? ( n63__$356 ) : ( cache_state ) ;
assign n65__$326 =  ( n60__$136 ) == ( 1'b1 )  ;
assign n66__$328 =  ( cache_state ) == ( bv_2_2_n10__$63 )  ;
assign n67__$330 = ~ ( n66__$328 )  ;
assign n68__$331 =  ( n67__$330 ) | ( n42__$124 )  ;
assign n69__$332 =  ( n65__$326 ) & (n68__$331 )  ;
assign n70__$333 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign n71__$335 = ~ ( n70__$333 )  ;
assign n72__$336 =  ( n69__$332 ) & (n71__$335 )  ;
assign n73__$366 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n74__$368 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n75__$370 =  ( n74__$368 ) ? ( msg1_source ) : ( cur_msg_source ) ;
assign n76__$371 =  ( n73__$366 ) ? ( n75__$370 ) : ( cache_owner ) ;
assign n77__$372 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign n79__$376 = nondet___unknown__1_n78 ;
assign n80__$392 =  ( n77__$372 ) ? ( n79__$376 ) : ( cache_owner ) ;
assign n81__$393 =  ( n72__$336 ) ? ( n76__$371 ) : ( n80__$392 ) ;
assign n82__$349 =  ( n72__$336 ) ? ( bv_2_0_n6__$59 ) : ( bv_2_1_n31__$97 ) ;
assign n83__$337 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n84__$339 =  ( n72__$336 ) | ( n83__$337 )  ;
assign n85__$340 =  ( n84__$339 ) ? ( cur_msg_type ) : ( msg1_type ) ;
assign n86__$345 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n87__$347 =  ( n72__$336 ) | ( n86__$345 )  ;
assign n88__$348 =  ( n87__$347 ) ? ( cur_msg_source ) : ( msg1_source ) ;
assign n89__$341 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n90__$343 =  ( n72__$336 ) | ( n89__$341 )  ;
assign n91__$344 =  ( n90__$343 ) ? ( cur_msg_tag ) : ( msg1_tag ) ;
always @(posedge clk) begin
   if(rst) begin
       msg1_ready <= msg1_ready_randinit ;
       msg3_ready <= msg3_ready_randinit ;
       msg2_type <= msg2_type_randinit ;
       msg2_valid <= msg2_valid_randinit ;
       cache_tag <= cache_tag_randinit ;
       cache_vd <= cache_vd_randinit ;
       cache_state <= cache_state_randinit ;
       cache_data <= cache_data_randinit ;
       cache_owner <= cache_owner_randinit ;
       share_list <= share_list_randinit ;
       cur_msg_state <= cur_msg_state_randinit ;
       cur_msg_type <= cur_msg_type_randinit ;
       cur_msg_source <= cur_msg_source_randinit ;
       cur_msg_tag <= cur_msg_tag_randinit ;
       __COUNTER_start__n15 <= 0;
   end
   else if(__START__ && __ILA_PMESH_L2_ILA_valid__) begin
       if ( __ILA_PMESH_L2_ILA_decode_of_STORE_REQ__ ) begin 
           __COUNTER_start__n15 <= 1; end
       else if( (__COUNTER_start__n15 >= 1 ) && ( __COUNTER_start__n15 < 255 )) begin
           __COUNTER_start__n15 <= __COUNTER_start__n15 + 1; end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           msg1_ready <= msg1_ready ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           msg3_ready <= msg3_ready ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           msg2_type <= n49__$419 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           msg2_valid <= msg2_valid ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cache_tag <= cache_tag ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cache_vd <= n53__$365 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cache_state <= n64__$357 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cache_data <= cache_data ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cache_owner <= n81__$393 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           share_list <= share_list ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cur_msg_state <= n82__$349 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cur_msg_type <= n85__$340 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cur_msg_source <= n88__$348 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_STORE_REQ__) begin
           cur_msg_tag <= n91__$344 ;
       end
   end
end
endmodule
