module PMESH_L2_ILA__DOT__LOAD_REQ(
__START__,
clk,
msg1_data,
msg1_source,
msg1_tag,
msg1_type,
msg1_valid,
msg2_ready,
msg3_data,
msg3_source,
msg3_tag,
msg3_type,
msg3_valid,
nondet___unknown__0_n76,
rst,
__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__,
__ILA_PMESH_L2_ILA_valid__,
msg1_ready,
msg3_ready,
msg2_type,
msg2_valid,
cache_tag,
cache_vd,
cache_state,
cache_data,
cache_owner,
share_list,
cur_msg_state,
cur_msg_type,
cur_msg_source,
cur_msg_tag,
__COUNTER_start__n15
);
input            __START__;
input            clk;
input     [63:0] msg1_data;
input      [5:0] msg1_source;
input     [25:0] msg1_tag;
input      [7:0] msg1_type;
input            msg1_valid;
input            msg2_ready;
input     [63:0] msg3_data;
input      [5:0] msg3_source;
input     [25:0] msg3_tag;
input      [7:0] msg3_type;
input            msg3_valid;
input      [5:0] nondet___unknown__0_n76;
input            rst;
output            __ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__;
output            __ILA_PMESH_L2_ILA_valid__;
output reg            msg1_ready;
output reg            msg3_ready;
output reg      [7:0] msg2_type;
output reg            msg2_valid;
output reg     [25:0] cache_tag;
output reg      [1:0] cache_vd;
output reg      [1:0] cache_state;
output reg     [63:0] cache_data;
output reg      [5:0] cache_owner;
output reg     [63:0] share_list;
output reg      [1:0] cur_msg_state;
output reg      [7:0] cur_msg_type;
output reg      [5:0] cur_msg_source;
output reg     [25:0] cur_msg_tag;
output reg      [7:0] __COUNTER_start__n15;
wire            __ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__;
wire            __ILA_PMESH_L2_ILA_valid__;
wire            __START__;
wire            bv_1_1_n0__$172;
wire      [1:0] bv_2_0_n6__$59;
wire      [1:0] bv_2_1_n31__$97;
wire      [1:0] bv_2_2_n10__$63;
wire      [1:0] bv_2_3_n21__$105;
wire     [63:0] bv_64_1_n82__$269;
wire      [7:0] bv_8_16_n44__$73;
wire      [7:0] bv_8_17_n34__$75;
wire      [7:0] bv_8_18_n33__$77;
wire      [7:0] bv_8_19_n29__$79;
wire      [7:0] bv_8_20_n28__$81;
wire      [7:0] bv_8_29_n43__$93;
wire      [7:0] bv_8_31_n4__$67;
(* keep *) wire     [63:0] cache_data_randinit;
(* keep *) wire      [5:0] cache_owner_randinit;
(* keep *) wire      [1:0] cache_state_randinit;
(* keep *) wire     [25:0] cache_tag_randinit;
(* keep *) wire      [1:0] cache_vd_randinit;
wire            clk;
(* keep *) wire      [5:0] cur_msg_source_randinit;
(* keep *) wire      [1:0] cur_msg_state_randinit;
(* keep *) wire     [25:0] cur_msg_tag_randinit;
(* keep *) wire      [7:0] cur_msg_type_randinit;
wire     [63:0] msg1_data;
(* keep *) wire            msg1_ready_randinit;
wire      [5:0] msg1_source;
wire     [25:0] msg1_tag;
wire      [7:0] msg1_type;
wire            msg1_valid;
wire            msg2_ready;
(* keep *) wire      [7:0] msg2_type_randinit;
(* keep *) wire            msg2_valid_randinit;
wire     [63:0] msg3_data;
(* keep *) wire            msg3_ready_randinit;
wire      [5:0] msg3_source;
wire     [25:0] msg3_tag;
wire      [7:0] msg3_type;
wire            msg3_valid;
wire            n11__$188;
wire            n12__$190;
wire            n13__$191;
wire            n14__$192;
wire            n16__$137;
wire     [25:0] n17__$139;
wire            n18__$140;
wire            n19__$142;
wire            n1__$174;
wire            n20__$143;
wire            n22__$145;
wire            n23__$147;
wire            n24__$148;
wire            n25__$281;
wire            n26__$283;
wire            n27__$285;
wire            n2__$178;
wire      [7:0] n30__$287;
wire            n32__$288;
wire      [7:0] n35__$290;
wire      [7:0] n36__$291;
wire            n37__$149;
wire            n38__$294;
wire            n39__$296;
wire            n3__$180;
wire            n40__$121;
wire      [5:0] n41__$123;
wire            n42__$124;
wire      [7:0] n45__$298;
wire      [7:0] n46__$299;
wire      [7:0] n47__$300;
wire      [7:0] n48__$301;
wire            n49__$260;
wire            n50__$262;
wire      [1:0] n51__$264;
wire      [1:0] n52__$265;
wire            n53__$126;
wire     [25:0] n54__$128;
wire            n55__$129;
wire            n56__$131;
wire            n57__$133;
wire            n58__$135;
wire            n59__$136;
wire            n5__$181;
wire            n60__$219;
wire            n61__$221;
wire      [1:0] n62__$223;
wire      [1:0] n63__$224;
wire            n64__$195;
wire            n65__$197;
wire            n66__$199;
wire            n67__$200;
wire            n68__$201;
wire            n69__$225;
wire            n70__$227;
wire      [5:0] n71__$229;
wire      [5:0] n72__$230;
wire            n73__$233;
wire            n74__$235;
wire            n75__$237;
wire      [5:0] n77__$240;
wire      [5:0] n78__$256;
wire      [5:0] n79__$257;
wire            n7__$183;
wire            n80__$266;
wire            n81__$268;
wire            n83__$271;
wire      [5:0] n84__$273;
wire     [63:0] n85__$274;
wire     [63:0] n86__$276;
wire     [63:0] n87__$277;
wire     [63:0] n88__$278;
wire      [1:0] n89__$216;
wire            n8__$185;
wire            n90__$204;
wire            n91__$206;
wire      [7:0] n92__$207;
wire            n93__$212;
wire            n94__$214;
wire      [5:0] n95__$215;
wire            n96__$208;
wire            n97__$210;
wire     [25:0] n98__$211;
wire            n9__$186;
wire      [5:0] nondet___unknown__0_n76;
wire            rst;
(* keep *) wire     [63:0] share_list_randinit;
assign __ILA_PMESH_L2_ILA_valid__ = 1'b1 ;
assign bv_1_1_n0__$172 = 1'h1 ;
assign n1__$174 =  ( msg1_ready ) == ( bv_1_1_n0__$172 )  ;
assign n2__$178 =  ( msg1_valid ) == ( bv_1_1_n0__$172 )  ;
assign n3__$180 =  ( n1__$174 ) & (n2__$178 )  ;
assign bv_8_31_n4__$67 = 8'h1f ;
assign n5__$181 =  ( msg1_type ) == ( bv_8_31_n4__$67 )  ;
assign bv_2_0_n6__$59 = 2'h0 ;
assign n7__$183 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n8__$185 =  ( n5__$181 ) & (n7__$183 )  ;
assign n9__$186 =  ( cur_msg_type ) == ( bv_8_31_n4__$67 )  ;
assign bv_2_2_n10__$63 = 2'h2 ;
assign n11__$188 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n12__$190 =  ( n9__$186 ) & (n11__$188 )  ;
assign n13__$191 =  ( n8__$185 ) | ( n12__$190 )  ;
assign n14__$192 =  ( n3__$180 ) & (n13__$191 )  ;
assign __ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__ = n14__$192 ;
assign n16__$137 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n17__$139 =  ( n16__$137 ) ? ( msg1_tag ) : ( cur_msg_tag ) ;
assign n18__$140 =  ( n17__$139 ) == ( cache_tag )  ;
assign n19__$142 = ~ ( n18__$140 )  ;
assign n20__$143 =  ( cache_vd ) == ( bv_2_2_n10__$63 )  ;
assign bv_2_3_n21__$105 = 2'h3 ;
assign n22__$145 =  ( cache_vd ) == ( bv_2_3_n21__$105 )  ;
assign n23__$147 =  ( n20__$143 ) | ( n22__$145 )  ;
assign n24__$148 =  ( n19__$142 ) & (n23__$147 )  ;
assign n25__$281 =  ( n24__$148 ) == ( 1'b1 )  ;
assign n26__$283 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n27__$285 =  ( cache_vd ) == ( bv_2_3_n21__$105 )  ;
assign bv_8_20_n28__$81 = 8'h14 ;
assign bv_8_19_n29__$79 = 8'h13 ;
assign n30__$287 =  ( n27__$285 ) ? ( bv_8_20_n28__$81 ) : ( bv_8_19_n29__$79 ) ;
assign bv_2_1_n31__$97 = 2'h1 ;
assign n32__$288 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign bv_8_18_n33__$77 = 8'h12 ;
assign bv_8_17_n34__$75 = 8'h11 ;
assign n35__$290 =  ( n32__$288 ) ? ( bv_8_18_n33__$77 ) : ( bv_8_17_n34__$75 ) ;
assign n36__$291 =  ( n26__$283 ) ? ( n30__$287 ) : ( n35__$290 ) ;
assign n37__$149 =  ( cache_vd ) == ( bv_2_0_n6__$59 )  ;
assign n38__$294 =  ( n37__$149 ) == ( 1'b1 )  ;
assign n39__$296 =  ( cache_state ) == ( bv_2_2_n10__$63 )  ;
assign n40__$121 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n41__$123 =  ( n40__$121 ) ? ( msg1_source ) : ( cur_msg_source ) ;
assign n42__$124 =  ( n41__$123 ) == ( cache_owner )  ;
assign bv_8_29_n43__$93 = 8'h1d ;
assign bv_8_16_n44__$73 = 8'h10 ;
assign n45__$298 =  ( n42__$124 ) ? ( bv_8_29_n43__$93 ) : ( bv_8_16_n44__$73 ) ;
assign n46__$299 =  ( n39__$296 ) ? ( n45__$298 ) : ( bv_8_29_n43__$93 ) ;
assign n47__$300 =  ( n38__$294 ) ? ( bv_8_19_n29__$79 ) : ( n46__$299 ) ;
assign n48__$301 =  ( n25__$281 ) ? ( n36__$291 ) : ( n47__$300 ) ;
assign n49__$260 =  ( n24__$148 ) == ( 1'b1 )  ;
assign n50__$262 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n51__$264 =  ( n50__$262 ) ? ( bv_2_0_n6__$59 ) : ( cache_vd ) ;
assign n52__$265 =  ( n49__$260 ) ? ( n51__$264 ) : ( cache_vd ) ;
assign n53__$126 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n54__$128 =  ( n53__$126 ) ? ( msg1_tag ) : ( cur_msg_tag ) ;
assign n55__$129 =  ( n54__$128 ) == ( cache_tag )  ;
assign n56__$131 =  ( cache_vd ) == ( bv_2_2_n10__$63 )  ;
assign n57__$133 =  ( cache_vd ) == ( bv_2_3_n21__$105 )  ;
assign n58__$135 =  ( n56__$131 ) | ( n57__$133 )  ;
assign n59__$136 =  ( n55__$129 ) & (n58__$135 )  ;
assign n60__$219 =  ( n59__$136 ) == ( 1'b1 )  ;
assign n61__$221 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n62__$223 =  ( n61__$221 ) ? ( bv_2_2_n10__$63 ) : ( cache_state ) ;
assign n63__$224 =  ( n60__$219 ) ? ( n62__$223 ) : ( cache_state ) ;
assign n64__$195 =  ( n59__$136 ) == ( 1'b1 )  ;
assign n65__$197 =  ( cache_state ) == ( bv_2_2_n10__$63 )  ;
assign n66__$199 = ~ ( n65__$197 )  ;
assign n67__$200 =  ( n66__$199 ) | ( n42__$124 )  ;
assign n68__$201 =  ( n64__$195 ) & (n67__$200 )  ;
assign n69__$225 =  ( cache_state ) == ( bv_2_0_n6__$59 )  ;
assign n70__$227 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n71__$229 =  ( n70__$227 ) ? ( msg1_source ) : ( cur_msg_source ) ;
assign n72__$230 =  ( n69__$225 ) ? ( n71__$229 ) : ( cache_owner ) ;
assign n73__$233 =  ( n24__$148 ) == ( 1'b1 )  ;
assign n74__$235 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign n75__$237 =  ( n73__$233 ) & (n74__$235 )  ;
assign n77__$240 = nondet___unknown__0_n76 ;
assign n78__$256 =  ( n75__$237 ) ? ( n77__$240 ) : ( cache_owner ) ;
assign n79__$257 =  ( n68__$201 ) ? ( n72__$230 ) : ( n78__$256 ) ;
assign n80__$266 =  ( cache_state ) == ( bv_2_1_n31__$97 )  ;
assign n81__$268 =  ( n68__$201 ) & (n80__$266 )  ;
assign bv_64_1_n82__$269 = 64'h1 ;
assign n83__$271 =  ( cur_msg_state ) == ( bv_2_0_n6__$59 )  ;
assign n84__$273 =  ( n83__$271 ) ? ( msg1_source ) : ( cur_msg_source ) ;
assign n85__$274 =  {58'd0 , n84__$273}  ;
assign n86__$276 =  ( bv_64_1_n82__$269 ) << ( n85__$274 )  ;
assign n87__$277 =  ( share_list ) | ( n86__$276 )  ;
assign n88__$278 =  ( n81__$268 ) ? ( n87__$277 ) : ( share_list ) ;
assign n89__$216 =  ( n68__$201 ) ? ( bv_2_0_n6__$59 ) : ( bv_2_1_n31__$97 ) ;
assign n90__$204 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n91__$206 =  ( n68__$201 ) | ( n90__$204 )  ;
assign n92__$207 =  ( n91__$206 ) ? ( cur_msg_type ) : ( msg1_type ) ;
assign n93__$212 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n94__$214 =  ( n68__$201 ) | ( n93__$212 )  ;
assign n95__$215 =  ( n94__$214 ) ? ( cur_msg_source ) : ( msg1_source ) ;
assign n96__$208 =  ( cur_msg_state ) == ( bv_2_2_n10__$63 )  ;
assign n97__$210 =  ( n68__$201 ) | ( n96__$208 )  ;
assign n98__$211 =  ( n97__$210 ) ? ( cur_msg_tag ) : ( msg1_tag ) ;
always @(posedge clk) begin
   if(rst) begin
       msg1_ready <= msg1_ready_randinit ;
       msg3_ready <= msg3_ready_randinit ;
       msg2_type <= msg2_type_randinit ;
       msg2_valid <= msg2_valid_randinit ;
       cache_tag <= cache_tag_randinit ;
       cache_vd <= cache_vd_randinit ;
       cache_state <= cache_state_randinit ;
       cache_data <= cache_data_randinit ;
       cache_owner <= cache_owner_randinit ;
       share_list <= share_list_randinit ;
       cur_msg_state <= cur_msg_state_randinit ;
       cur_msg_type <= cur_msg_type_randinit ;
       cur_msg_source <= cur_msg_source_randinit ;
       cur_msg_tag <= cur_msg_tag_randinit ;
       __COUNTER_start__n15 <= 0;
   end
   else if(__START__ && __ILA_PMESH_L2_ILA_valid__) begin
       if ( __ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__ ) begin 
           __COUNTER_start__n15 <= 1; end
       else if( (__COUNTER_start__n15 >= 1 ) && ( __COUNTER_start__n15 < 255 )) begin
           __COUNTER_start__n15 <= __COUNTER_start__n15 + 1; end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           msg1_ready <= msg1_ready ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           msg3_ready <= msg3_ready ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           msg2_type <= n48__$301 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           msg2_valid <= bv_1_1_n0__$172 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cache_tag <= cache_tag ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cache_vd <= n52__$265 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cache_state <= n63__$224 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cache_data <= cache_data ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cache_owner <= n79__$257 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           share_list <= n88__$278 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cur_msg_state <= n89__$216 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cur_msg_type <= n92__$207 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cur_msg_source <= n95__$215 ;
       end
       if (__ILA_PMESH_L2_ILA_decode_of_LOAD_REQ__) begin
           cur_msg_tag <= n98__$211 ;
       end
   end
end
endmodule
